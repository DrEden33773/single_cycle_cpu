module mips (
    clk,
    rst
);

  input clk;  // clock
  input rst;  // reset

endmodule
